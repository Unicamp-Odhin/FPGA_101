module top (
    input  logic clk,  // 100MHz
    output logic [15:0] LED,
    input  logic [15:0] SW,
    input  logic CPU_RESETN
);



endmodule

