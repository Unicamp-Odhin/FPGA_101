module top (
    input logic clk,  // board clock 25mhz 

    output logic [7:0] LED
);

endmodule

